module usv_tb; 

	reg s1;
    reg s0;
    reg clk;
	reg [63:0]d;
    wire [63:0]q; 