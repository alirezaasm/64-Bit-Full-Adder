module ram (Data,
            address,
            data_out
            );
		
    parameter address_size = 64;
    parameter data_size    = 32;
	
	 input reg [address_size-1:0] Data [data_size-1 : 0];


endmodule