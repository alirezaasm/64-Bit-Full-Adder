module ram (Data,
            address,
            data_out
            );


endmodule