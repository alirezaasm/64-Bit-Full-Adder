module ram (Data,
            address

            );


endmodule