module FullAdder1 (
    input A,
    input B,
    input Cin,//input carry 
    output S,// sum 
    output Cout//out carry
	
	
    );

   

endmodule