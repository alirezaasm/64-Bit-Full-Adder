module usv_tb; 