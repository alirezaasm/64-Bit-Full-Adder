module ram (Data,
            address,
            data_out
            );
		
    parameter address_size = 64;
    parameter data_size    = 32;


endmodule