`include "./ram.v"
`include "../counter/Counter.v"

module ram_tb;
		
	reg clk, reset,s[1:0], data_in, SISR, SISL,
    reg reg_data;







endmodule
