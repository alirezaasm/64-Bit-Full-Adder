module usv_tb; 

	reg s1;
    reg s0;
    reg clk;