module ram (Data,
            );


endmodule