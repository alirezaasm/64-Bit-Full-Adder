module usv_tb;
